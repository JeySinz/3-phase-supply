CircuitMaker Text
5.6
Probes: 3
V1_1
Transient Analysis
0 445 200 65280
V3_1
Transient Analysis
1 564 204 65535
V4_1
Transient Analysis
2 664 224 16776960
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
270 120 30 100 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.419790 0.500000
344 176 1532 456
9961490 0
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 479 427 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7361 0 0
2
45139.4 0
0
11 Signal Gen~
195 354 373 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1012557331 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 250 0.01333 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V4
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 13.33m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
4747 0 0
2
45139.4 0
0
11 Signal Gen~
195 354 288 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
1004170870 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 250 0.006666 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
43 %D %1 %2 DC 0 SIN(0 250 50 6.666m 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
45139.4 0
0
11 Signal Gen~
195 352 205 0 19 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1132068864
20
1 50 0 250 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -250/250V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 250 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3472 0 0
2
45139.4 0
0
9 Resistor~
219 695 183 0 4 5
0 5 2 0 -1
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9998 0 0
2
45139.4 0
0
9 Resistor~
219 592 187 0 4 5
0 4 2 0 -1
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3536 0 0
2
45139.4 0
0
9 Resistor~
219 507 188 0 2 5
0 3 6
0
0 0 880 0
4 100k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 512 0 0 0 0
1 R
4597 0 0
2
45139.4 0
0
9
2 0 2 0 0 8192 0 3 0 0 3 4
385 293
444 293
444 390
479 390
2 0 2 0 0 8192 0 4 0 0 3 4
383 210
412 210
412 399
479 399
0 0 2 0 0 0 0 0 0 0 4 4
528 189
528 247
479 247
479 401
2 0 2 0 0 4096 0 6 0 0 5 5
610 187
610 390
471 390
471 401
479 401
2 0 2 0 0 12416 0 5 0 0 9 4
713 183
732 183
732 401
479 401
1 1 3 0 0 4224 0 4 7 0 0 4
383 200
467 200
467 188
489 188
1 1 4 0 0 4224 0 3 6 0 0 4
385 283
565 283
565 187
574 187
1 1 5 0 0 4224 0 2 5 0 0 4
385 368
665 368
665 183
677 183
2 1 2 0 0 0 0 2 1 0 0 3
385 378
479 378
479 421
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
